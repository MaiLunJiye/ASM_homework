module multi8 (in1, in2, out);
input reg[7:0] in1,in2;
output reg[15:0] out;
parameter lenth = 7;    //8 位长度

always @ (in1, in2)
begin

end

endmodule
