module mov(clk50hz, sw0, hex0, hex1, hex2);//input clk1hz,sw0;parameters Value=55'b0001001_0110000_1110001_1110001_0000001_0000000_0000000_0000000;//HELLO___output [6:0] hex0,hex1,hex2;reg[55:0] m=Valuealways @ (posedoge clk50hz)begin if (sw0) m = {m,m[55:49]}; else  m = {m[6:0],m[55:7]}; {hex0,hex1,hex2} = m[55:35];endendmodulemodule dicCLK(clk50,clk1);input clk50;output clk1;integer i;reg clk1;reg cs;always @ (posdege clk50)begin if (i==59) begin i=0; else i=i+1; if(i==59)endendmodule
