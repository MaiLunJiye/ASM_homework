module displayLed(num, outcode);
    input reg[3:0] num;
    output reg[6:0] outcode;

    always @ (num)
    begin
        case(num)
            4'b000: num=
    end
endmodule
